library verilog;
use verilog.vl_types.all;
entity Subsistema_4_vlg_vec_tst is
end Subsistema_4_vlg_vec_tst;
