library verilog;
use verilog.vl_types.all;
entity paralelo_serie_384b_vlg_check_tst is
    port(
        serial_out      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end paralelo_serie_384b_vlg_check_tst;
