library verilog;
use verilog.vl_types.all;
entity paralelo_serie_384b_vlg_vec_tst is
end paralelo_serie_384b_vlg_vec_tst;
