-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Mon Nov 10 16:18:45 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY subsistema2esquematico IS 
	PORT
	(
		inclk0 :  IN  STD_LOGIC;
		areset :  IN  STD_LOGIC;
		INICIO :  IN  STD_LOGIC;
		MV :  IN  STD_LOGIC;
		MINV :  IN  STD_LOGIC;
		TURNO :  IN  STD_LOGIC;
		VF :  IN  STD_LOGIC;
		VICTORIA :  IN  STD_LOGIC;
		EMPATE :  IN  STD_LOGIC;
		POSICION :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		SC1 :  IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
		SC2 :  IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
		CERO :  OUT  STD_LOGIC;
		UNO :  OUT  STD_LOGIC;
		locked :  OUT  STD_LOGIC;
		Y :  OUT  STD_LOGIC
	);
END subsistema2esquematico;

ARCHITECTURE bdf_type OF subsistema2esquematico IS 

COMPONENT block1
	PORT(inclk0 : IN STD_LOGIC;
		 areset : IN STD_LOGIC;
		 load : IN STD_LOGIC;
		 parallel_in : IN STD_LOGIC_VECTOR(383 DOWNTO 0);
		 CERO : OUT STD_LOGIC;
		 UNO : OUT STD_LOGIC;
		 frecuencialed : OUT STD_LOGIC;
		 locked : OUT STD_LOGIC;
		 Y : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT coloress2
	PORT(INICIO : IN STD_LOGIC;
		 MV : IN STD_LOGIC;
		 MINV : IN STD_LOGIC;
		 TURNO : IN STD_LOGIC;
		 VF : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 VICTORIA : IN STD_LOGIC;
		 EMPATE : IN STD_LOGIC;
		 POSICION : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 SC1 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 SC2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 MATRIZ : OUT STD_LOGIC_VECTOR(383 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_counter0
	PORT(clock : IN STD_LOGIC;
		 cout : OUT STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(383 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;


BEGIN 



b2v_inst : block1
PORT MAP(inclk0 => inclk0,
		 areset => areset,
		 load => SYNTHESIZED_WIRE_0,
		 parallel_in => SYNTHESIZED_WIRE_1,
		 CERO => CERO,
		 UNO => UNO,
		 frecuencialed => SYNTHESIZED_WIRE_4,
		 locked => locked,
		 Y => Y);


b2v_inst1 : coloress2
PORT MAP(INICIO => INICIO,
		 MV => MV,
		 MINV => MINV,
		 TURNO => TURNO,
		 VF => VF,
		 CLK => SYNTHESIZED_WIRE_4,
		 VICTORIA => VICTORIA,
		 EMPATE => EMPATE,
		 POSICION => POSICION,
		 SC1 => SC1,
		 SC2 => SC2,
		 MATRIZ => SYNTHESIZED_WIRE_1);


b2v_inst2 : lpm_counter0
PORT MAP(clock => SYNTHESIZED_WIRE_4,
		 cout => SYNTHESIZED_WIRE_0);


END bdf_type;