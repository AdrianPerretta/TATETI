library verilog;
use verilog.vl_types.all;
entity Detector_Victoria_vlg_vec_tst is
end Detector_Victoria_vlg_vec_tst;
