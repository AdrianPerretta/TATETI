library verilog;
use verilog.vl_types.all;
entity Validar_movimiento_vlg_vec_tst is
end Validar_movimiento_vlg_vec_tst;
