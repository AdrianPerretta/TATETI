library verilog;
use verilog.vl_types.all;
entity Colores_vlg_vec_tst is
end Colores_vlg_vec_tst;
