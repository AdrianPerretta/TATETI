library verilog;
use verilog.vl_types.all;
entity teclado_vlg_vec_tst is
end teclado_vlg_vec_tst;
